`include "master.sv"
`include "slave.sv"

module Master_AXI3 (
    input logic clk, rst,
    
);
    
Master 

endmodule